`ifndef I2C_IF_INCLUDED_
`define I2C_IF_INCLUDED_
//--------------------------------------------------------------------------------------------
// class     : I2C_intf
// Description  : Declaring the signals for i2c interface
//--------------------------------------------------------------------------------------------
interface i2c_if;


/*logic scl;
  logic sda;
  logic scl_i;
  logic sda_i;
 */

endinterface : i2c_if

`endif
